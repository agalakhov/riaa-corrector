.MODEL Swx ASWITCH(RON=1 ROFF=1 VON=1 VOFF=1)
R1 0 1 1MEG
AS1 0 1 2 3 Swx
R2 1 2 1MEG
R3 2 3 1MEG
R4 3 0 1MEG
